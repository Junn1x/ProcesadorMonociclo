module IM (
    input logic [31:0] address,
    output logic [31:0] inst
);

endmodule

