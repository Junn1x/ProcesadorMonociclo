module DM (
    input logic [31:0] address,
    input logic [31:0] DataWr,
    input logic DmWr,
    input logic [2:0] DmCtrl,
    output logic [31:0] DataRd
);

endmodule