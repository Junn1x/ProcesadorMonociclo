module PC (
    input logic [31:0] nextPcAdress,
    input logic clk,
    output logic [31:0] address
);


endmodule
